module main

// do.v -> Undo & Redo
struct Change {
}

fn describe_change() {
}

fn undo() {
}

fn redo() {
}
