module main

fn em_open_dialog() {
}
